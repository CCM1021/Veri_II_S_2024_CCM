package router_env_pkg;
import uvm_pkg::*;
import router_stimulus_pkg::*;
`include "labs\lab2\driver.sv"
`include "labs\lab2\input_agent.sv"
`include "labs\lab2\router_env.sv"
endpackage
